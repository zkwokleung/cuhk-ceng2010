library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity d2_counter_tb is
--  Port ( );
end d2_counter_tb;

architecture Behavioral of d2_counter_tb is

begin


end Behavioral;
